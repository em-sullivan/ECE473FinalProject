module controller (

	input [31:0] ins,
	output reg reg_wen,
	output reg reg_des,
	output reg jr,
	output reg [3:0] alu_code);
	
	
	always @* begin

	end
	
endmodule
